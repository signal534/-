module q1 (
    input [31:0] data_in,
    output reg [5:0] data_out
  );

  always @(*)
  begin
    casez (data_in)
      32'b1??????????????????????????????? :
        data_out = 6'd0;
      32'b01?????????????????????????????? :
        data_out = 6'd1;
      32'b001????????????????????????????? :
        data_out = 6'd2;
      32'b0001???????????????????????????? :
        data_out = 6'd3;
      32'b00001??????????????????????????? :
        data_out = 6'd4;
      32'b000001?????????????????????????? :
        data_out = 6'd5;
      32'b0000001????????????????????????? :
        data_out = 6'd6;
      32'b00000001???????????????????????? :
        data_out = 6'd7;
      32'b000000001??????????????????????? :
        data_out = 6'd8;
      32'b0000000001?????????????????????? :
        data_out = 6'd9;
      32'b00000000001????????????????????? :
        data_out = 6'd10;
      32'b000000000001???????????????????? :
        data_out = 6'd11;
      32'b0000000000001??????????????????? :
        data_out = 6'd12;
      32'b00000000000001?????????????????? :
        data_out = 6'd13;
      32'b000000000000001????????????????? :
        data_out = 6'd14;
      32'b0000000000000001???????????????? :
        data_out = 6'd15;
      32'b00000000000000001??????????????? :
        data_out = 6'd16;
      32'b000000000000000001?????????????? :
        data_out = 6'd17;
      32'b0000000000000000001????????????? :
        data_out = 6'd18;
      32'b00000000000000000001???????????? :
        data_out = 6'd19;
      32'b000000000000000000001??????????? :
        data_out = 6'd20;
      32'b0000000000000000000001?????????? :
        data_out = 6'd21;
      32'b00000000000000000000001????????? :
        data_out = 6'd22;
      32'b000000000000000000000001???????? :
        data_out = 6'd23;
      32'b0000000000000000000000001??????? :
        data_out = 6'd24;
      32'b00000000000000000000000001?????? :
        data_out = 6'd25;
      32'b000000000000000000000000001????? :
        data_out = 6'd26;
      32'b0000000000000000000000000001???? :
        data_out = 6'd27;
      32'b00000000000000000000000000001??? :
        data_out = 6'd28;
      32'b000000000000000000000000000001?? :
        data_out = 6'd29;
      32'b0000000000000000000000000000001? :
        data_out = 6'd30;
      32'b00000000000000000000000000000001 :
        data_out = 6'd31;
      default :
        data_out = 6'd32;
    endcase
  end

endmodule
